// system_0.v

// Generated using ACDS version 11.1sp2 259 at 2012.10.15.16:11:46

`timescale 1 ps / 1 ps
module system_0 (
		inout  wire [15:0] sram_16bit_512k_0_avalon_slave_0_export_DQ,                  // sram_16bit_512k_0_avalon_slave_0_export.DQ
		output wire [17:0] sram_16bit_512k_0_avalon_slave_0_export_ADDR,                //                                        .ADDR
		output wire        sram_16bit_512k_0_avalon_slave_0_export_UB_N,                //                                        .UB_N
		output wire        sram_16bit_512k_0_avalon_slave_0_export_LB_N,                //                                        .LB_N
		output wire        sram_16bit_512k_0_avalon_slave_0_export_WE_N,                //                                        .WE_N
		output wire        sram_16bit_512k_0_avalon_slave_0_export_CE_N,                //                                        .CE_N
		output wire        sram_16bit_512k_0_avalon_slave_0_export_OE_N,                //                                        .OE_N
		input  wire        clk_clk_in_reset_reset_n,                                    //                        clk_clk_in_reset.reset_n
		output wire        sd_clk_external_connection_export,                           //              sd_clk_external_connection.export
		output wire [9:0]  led_red_external_connection_export,                          //             led_red_external_connection.export
		inout  wire        sd_dat_external_connection_export,                           //              sd_dat_external_connection.export
		output wire [11:0] sdram_0_wire_addr,                                           //                            sdram_0_wire.addr
		output wire [1:0]  sdram_0_wire_ba,                                             //                                        .ba
		output wire        sdram_0_wire_cas_n,                                          //                                        .cas_n
		output wire        sdram_0_wire_cke,                                            //                                        .cke
		output wire        sdram_0_wire_cs_n,                                           //                                        .cs_n
		inout  wire [15:0] sdram_0_wire_dq,                                             //                                        .dq
		output wire [1:0]  sdram_0_wire_dqm,                                            //                                        .dqm
		output wire        sdram_0_wire_ras_n,                                          //                                        .ras_n
		output wire        sdram_0_wire_we_n,                                           //                                        .we_n
		output wire [6:0]  seg7_display_conduit_end_oSEG0,                              //                seg7_display_conduit_end.oSEG0
		output wire [6:0]  seg7_display_conduit_end_oSEG1,                              //                                        .oSEG1
		output wire [6:0]  seg7_display_conduit_end_oSEG2,                              //                                        .oSEG2
		output wire [6:0]  seg7_display_conduit_end_oSEG3,                              //                                        .oSEG3
		output wire [6:0]  seg7_display_conduit_end_oSEG4,                              //                                        .oSEG4
		output wire [6:0]  seg7_display_conduit_end_oSEG5,                              //                                        .oSEG5
		output wire [6:0]  seg7_display_conduit_end_oSEG6,                              //                                        .oSEG6
		output wire [6:0]  seg7_display_conduit_end_oSEG7,                              //                                        .oSEG7
		inout  wire [7:0]  tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data,     //         tri_state_bridge_0_bridge_0_out.tri_state_bridge_0_data
		output wire        tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn,    //                                        .tri_state_bridge_0_readn
		output wire        tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0,  //                                        .write_n_to_the_cfi_flash_0
		output wire [21:0] tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address,  //                                        .tri_state_bridge_0_address
		output wire        tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0, //                                        .select_n_to_the_cfi_flash_0
		input  wire [3:0]  button_pio_external_connection_export,                       //          button_pio_external_connection.export
		output wire [7:0]  led_green_external_connection_export,                        //           led_green_external_connection.export
		input  wire        clk_clk_in_clk,                                              //                              clk_clk_in.clk
		output wire        audio_0_avalon_slave_0_export_oAUD_DATA,                     //           audio_0_avalon_slave_0_export.oAUD_DATA
		output wire        audio_0_avalon_slave_0_export_oAUD_LRCK,                     //                                        .oAUD_LRCK
		output wire        audio_0_avalon_slave_0_export_oAUD_BCK,                      //                                        .oAUD_BCK
		output wire        audio_0_avalon_slave_0_export_oAUD_XCK,                      //                                        .oAUD_XCK
		input  wire        audio_0_avalon_slave_0_export_iCLK_18_4,                     //                                        .iCLK_18_4
		input  wire [17:0] switch_pio_external_connection_export,                       //          switch_pio_external_connection.export
		input  wire        uart_0_external_connection_rxd,                              //              uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd,                              //                                        .txd
		inout  wire        sd_cmd_external_connection_export                            //              sd_cmd_external_connection.export
	);

	wire   [0:0] tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out;                                     // tri_state_bridge_0_pinSharer_0:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0:tcs_select_n_to_the_cfi_flash_0
	wire  [21:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out;                                      // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_address -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_address
	wire         tri_state_bridge_0_pinsharer_0_tcm_grant;                                                               // tri_state_bridge_0_bridge_0:grant -> tri_state_bridge_0_pinSharer_0:grant
	wire   [0:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out;                                        // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_readn -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_readn
	wire         tri_state_bridge_0_pinsharer_0_tcm_request;                                                             // tri_state_bridge_0_pinSharer_0:request -> tri_state_bridge_0_bridge_0:request
	wire   [7:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in;                                          // tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data_in -> tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data_in
	wire         tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen;                                       // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data_outen -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data_outen
	wire   [0:0] tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out;                                      // tri_state_bridge_0_pinSharer_0:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0:tcs_write_n_to_the_cfi_flash_0
	wire   [7:0] tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out;                                         // tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data
	wire         cfi_flash_0_tcm_chipselect_n_out;                                                                       // cfi_flash_0:tcm_chipselect_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_chipselect_n_out
	wire         cfi_flash_0_tcm_grant;                                                                                  // tri_state_bridge_0_pinSharer_0:tcs0_grant -> cfi_flash_0:tcm_grant
	wire         cfi_flash_0_tcm_data_outen;                                                                             // cfi_flash_0:tcm_data_outen -> tri_state_bridge_0_pinSharer_0:tcs0_data_outen
	wire         cfi_flash_0_tcm_request;                                                                                // cfi_flash_0:tcm_request -> tri_state_bridge_0_pinSharer_0:tcs0_request
	wire   [7:0] cfi_flash_0_tcm_data_out;                                                                               // cfi_flash_0:tcm_data_out -> tri_state_bridge_0_pinSharer_0:tcs0_data_out
	wire         cfi_flash_0_tcm_write_n_out;                                                                            // cfi_flash_0:tcm_write_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_write_n_out
	wire  [21:0] cfi_flash_0_tcm_address_out;                                                                            // cfi_flash_0:tcm_address_out -> tri_state_bridge_0_pinSharer_0:tcs0_address_out
	wire   [7:0] cfi_flash_0_tcm_data_in;                                                                                // tri_state_bridge_0_pinSharer_0:tcs0_data_in -> cfi_flash_0:tcm_data_in
	wire         cfi_flash_0_tcm_read_n_out;                                                                             // cfi_flash_0:tcm_read_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_read_n_out
	wire         nios2_qsys_0_instruction_master_waitrequest;                                                            // nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [24:0] nios2_qsys_0_instruction_master_address;                                                                // nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	wire         nios2_qsys_0_instruction_master_read;                                                                   // nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                                               // nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_readdatavalid;                                                          // nios2_qsys_0_instruction_master_translator:av_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire         nios2_qsys_0_data_master_waitrequest;                                                                   // nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                                                     // nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	wire  [24:0] nios2_qsys_0_data_master_address;                                                                       // nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	wire         nios2_qsys_0_data_master_write;                                                                         // nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	wire         nios2_qsys_0_data_master_read;                                                                          // nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                                                      // nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                                                                   // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	wire         nios2_qsys_0_data_master_readdatavalid;                                                                 // nios2_qsys_0_data_master_translator:av_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                                                    // nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                // nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                  // nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                               // nios2_qsys_0_jtag_debug_module_translator:av_chipselect -> nios2_qsys_0:jtag_debug_module_select
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                    // nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                 // nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                            // nios2_qsys_0_jtag_debug_module_translator:av_begintransfer -> nios2_qsys_0:jtag_debug_module_begintransfer
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                              // nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                               // nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire  [15:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                              // sram_16bit_512k_0_avalon_slave_0_translator:av_writedata -> sram_16bit_512k_0:iDATA
	wire  [17:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                // sram_16bit_512k_0_avalon_slave_0_translator:av_address -> sram_16bit_512k_0:iADDR
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                             // sram_16bit_512k_0_avalon_slave_0_translator:av_chipselect -> sram_16bit_512k_0:iCE_N
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                  // sram_16bit_512k_0_avalon_slave_0_translator:av_write -> sram_16bit_512k_0:iWE_N
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                   // sram_16bit_512k_0_avalon_slave_0_translator:av_read -> sram_16bit_512k_0:iOE_N
	wire  [15:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                               // sram_16bit_512k_0:oDATA -> sram_16bit_512k_0_avalon_slave_0_translator:av_readdata
	wire   [1:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                             // sram_16bit_512k_0_avalon_slave_0_translator:av_byteenable -> sram_16bit_512k_0:iBE_N
	wire  [31:0] epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata;                             // epcs_controller_epcs_control_port_translator:av_writedata -> epcs_controller:writedata
	wire   [8:0] epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address;                               // epcs_controller_epcs_control_port_translator:av_address -> epcs_controller:address
	wire         epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect;                            // epcs_controller_epcs_control_port_translator:av_chipselect -> epcs_controller:chipselect
	wire         epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write;                                 // epcs_controller_epcs_control_port_translator:av_write -> epcs_controller:write_n
	wire         epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read;                                  // epcs_controller_epcs_control_port_translator:av_read -> epcs_controller:read_n
	wire  [31:0] epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata;                              // epcs_controller:readdata -> epcs_controller_epcs_control_port_translator:av_readdata
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest;                                             // cfi_flash_0:uas_waitrequest -> cfi_flash_0_uas_translator:av_waitrequest
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount;                                              // cfi_flash_0_uas_translator:av_burstcount -> cfi_flash_0:uas_burstcount
	wire   [7:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata;                                               // cfi_flash_0_uas_translator:av_writedata -> cfi_flash_0:uas_writedata
	wire  [21:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_address;                                                 // cfi_flash_0_uas_translator:av_address -> cfi_flash_0:uas_address
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_lock;                                                    // cfi_flash_0_uas_translator:av_lock -> cfi_flash_0:uas_lock
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_write;                                                   // cfi_flash_0_uas_translator:av_write -> cfi_flash_0:uas_write
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_read;                                                    // cfi_flash_0_uas_translator:av_read -> cfi_flash_0:uas_read
	wire   [7:0] cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata;                                                // cfi_flash_0:uas_readdata -> cfi_flash_0_uas_translator:av_readdata
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess;                                             // cfi_flash_0_uas_translator:av_debugaccess -> cfi_flash_0:uas_debugaccess
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid;                                           // cfi_flash_0:uas_readdatavalid -> cfi_flash_0_uas_translator:av_readdatavalid
	wire         cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable;                                              // cfi_flash_0_uas_translator:av_byteenable -> cfi_flash_0:uas_byteenable
	wire         sdram_0_s1_translator_avalon_anti_slave_0_waitrequest;                                                  // sdram_0:za_waitrequest -> sdram_0_s1_translator:av_waitrequest
	wire  [15:0] sdram_0_s1_translator_avalon_anti_slave_0_writedata;                                                    // sdram_0_s1_translator:av_writedata -> sdram_0:az_data
	wire  [21:0] sdram_0_s1_translator_avalon_anti_slave_0_address;                                                      // sdram_0_s1_translator:av_address -> sdram_0:az_addr
	wire         sdram_0_s1_translator_avalon_anti_slave_0_chipselect;                                                   // sdram_0_s1_translator:av_chipselect -> sdram_0:az_cs
	wire         sdram_0_s1_translator_avalon_anti_slave_0_write;                                                        // sdram_0_s1_translator:av_write -> sdram_0:az_wr_n
	wire         sdram_0_s1_translator_avalon_anti_slave_0_read;                                                         // sdram_0_s1_translator:av_read -> sdram_0:az_rd_n
	wire  [15:0] sdram_0_s1_translator_avalon_anti_slave_0_readdata;                                                     // sdram_0:za_data -> sdram_0_s1_translator:av_readdata
	wire         sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid;                                                // sdram_0:za_valid -> sdram_0_s1_translator:av_readdatavalid
	wire   [1:0] sdram_0_s1_translator_avalon_anti_slave_0_byteenable;                                                   // sdram_0_s1_translator:av_byteenable -> sdram_0:az_be_n
	wire  [15:0] audio_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                        // Audio_0_avalon_slave_0_translator:av_writedata -> Audio_0:iDATA
	wire         audio_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                            // Audio_0_avalon_slave_0_translator:av_write -> Audio_0:iWR
	wire  [15:0] audio_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                         // Audio_0:oDATA -> Audio_0_avalon_slave_0_translator:av_readdata
	wire  [31:0] seg7_display_avalon_slave_translator_avalon_anti_slave_0_writedata;                                     // SEG7_Display_avalon_slave_translator:av_writedata -> SEG7_Display:iDIG
	wire         seg7_display_avalon_slave_translator_avalon_anti_slave_0_write;                                         // SEG7_Display_avalon_slave_translator:av_write -> SEG7_Display:iWR
	wire  [31:0] led_green_s1_translator_avalon_anti_slave_0_writedata;                                                  // led_green_s1_translator:av_writedata -> led_green:writedata
	wire   [1:0] led_green_s1_translator_avalon_anti_slave_0_address;                                                    // led_green_s1_translator:av_address -> led_green:address
	wire         led_green_s1_translator_avalon_anti_slave_0_chipselect;                                                 // led_green_s1_translator:av_chipselect -> led_green:chipselect
	wire         led_green_s1_translator_avalon_anti_slave_0_write;                                                      // led_green_s1_translator:av_write -> led_green:write_n
	wire  [31:0] led_green_s1_translator_avalon_anti_slave_0_readdata;                                                   // led_green:readdata -> led_green_s1_translator:av_readdata
	wire  [31:0] led_red_s1_translator_avalon_anti_slave_0_writedata;                                                    // led_red_s1_translator:av_writedata -> led_red:writedata
	wire   [1:0] led_red_s1_translator_avalon_anti_slave_0_address;                                                      // led_red_s1_translator:av_address -> led_red:address
	wire         led_red_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led_red_s1_translator:av_chipselect -> led_red:chipselect
	wire         led_red_s1_translator_avalon_anti_slave_0_write;                                                        // led_red_s1_translator:av_write -> led_red:write_n
	wire  [31:0] led_red_s1_translator_avalon_anti_slave_0_readdata;                                                     // led_red:readdata -> led_red_s1_translator:av_readdata
	wire  [31:0] sd_clk_s1_translator_avalon_anti_slave_0_writedata;                                                     // SD_CLK_s1_translator:av_writedata -> SD_CLK:writedata
	wire   [1:0] sd_clk_s1_translator_avalon_anti_slave_0_address;                                                       // SD_CLK_s1_translator:av_address -> SD_CLK:address
	wire         sd_clk_s1_translator_avalon_anti_slave_0_chipselect;                                                    // SD_CLK_s1_translator:av_chipselect -> SD_CLK:chipselect
	wire         sd_clk_s1_translator_avalon_anti_slave_0_write;                                                         // SD_CLK_s1_translator:av_write -> SD_CLK:write_n
	wire  [31:0] sd_clk_s1_translator_avalon_anti_slave_0_readdata;                                                      // SD_CLK:readdata -> SD_CLK_s1_translator:av_readdata
	wire  [31:0] sd_cmd_s1_translator_avalon_anti_slave_0_writedata;                                                     // SD_CMD_s1_translator:av_writedata -> SD_CMD:writedata
	wire   [1:0] sd_cmd_s1_translator_avalon_anti_slave_0_address;                                                       // SD_CMD_s1_translator:av_address -> SD_CMD:address
	wire         sd_cmd_s1_translator_avalon_anti_slave_0_chipselect;                                                    // SD_CMD_s1_translator:av_chipselect -> SD_CMD:chipselect
	wire         sd_cmd_s1_translator_avalon_anti_slave_0_write;                                                         // SD_CMD_s1_translator:av_write -> SD_CMD:write_n
	wire  [31:0] sd_cmd_s1_translator_avalon_anti_slave_0_readdata;                                                      // SD_CMD:readdata -> SD_CMD_s1_translator:av_readdata
	wire  [31:0] sd_dat_s1_translator_avalon_anti_slave_0_writedata;                                                     // SD_DAT_s1_translator:av_writedata -> SD_DAT:writedata
	wire   [1:0] sd_dat_s1_translator_avalon_anti_slave_0_address;                                                       // SD_DAT_s1_translator:av_address -> SD_DAT:address
	wire         sd_dat_s1_translator_avalon_anti_slave_0_chipselect;                                                    // SD_DAT_s1_translator:av_chipselect -> SD_DAT:chipselect
	wire         sd_dat_s1_translator_avalon_anti_slave_0_write;                                                         // SD_DAT_s1_translator:av_write -> SD_DAT:write_n
	wire  [31:0] sd_dat_s1_translator_avalon_anti_slave_0_readdata;                                                      // SD_DAT:readdata -> SD_DAT_s1_translator:av_readdata
	wire   [1:0] switch_pio_s1_translator_avalon_anti_slave_0_address;                                                   // switch_pio_s1_translator:av_address -> switch_pio:address
	wire  [31:0] switch_pio_s1_translator_avalon_anti_slave_0_readdata;                                                  // switch_pio:readdata -> switch_pio_s1_translator:av_readdata
	wire  [31:0] button_pio_s1_translator_avalon_anti_slave_0_writedata;                                                 // button_pio_s1_translator:av_writedata -> button_pio:writedata
	wire   [1:0] button_pio_s1_translator_avalon_anti_slave_0_address;                                                   // button_pio_s1_translator:av_address -> button_pio:address
	wire         button_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                // button_pio_s1_translator:av_chipselect -> button_pio:chipselect
	wire         button_pio_s1_translator_avalon_anti_slave_0_write;                                                     // button_pio_s1_translator:av_write -> button_pio:write_n
	wire  [31:0] button_pio_s1_translator_avalon_anti_slave_0_readdata;                                                  // button_pio:readdata -> button_pio_s1_translator:av_readdata
	wire  [15:0] timer_1_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_1_s1_translator:av_writedata -> timer_1:writedata
	wire   [2:0] timer_1_s1_translator_avalon_anti_slave_0_address;                                                      // timer_1_s1_translator:av_address -> timer_1:address
	wire         timer_1_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	wire         timer_1_s1_translator_avalon_anti_slave_0_write;                                                        // timer_1_s1_translator:av_write -> timer_1:write_n
	wire  [15:0] timer_1_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_1:readdata -> timer_1_s1_translator:av_readdata
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                    // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                      // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                   // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                        // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                     // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire  [15:0] uart_0_s1_translator_avalon_anti_slave_0_writedata;                                                     // uart_0_s1_translator:av_writedata -> uart_0:writedata
	wire   [2:0] uart_0_s1_translator_avalon_anti_slave_0_address;                                                       // uart_0_s1_translator:av_address -> uart_0:address
	wire         uart_0_s1_translator_avalon_anti_slave_0_chipselect;                                                    // uart_0_s1_translator:av_chipselect -> uart_0:chipselect
	wire         uart_0_s1_translator_avalon_anti_slave_0_write;                                                         // uart_0_s1_translator:av_write -> uart_0:write_n
	wire         uart_0_s1_translator_avalon_anti_slave_0_read;                                                          // uart_0_s1_translator:av_read -> uart_0:read_n
	wire  [15:0] uart_0_s1_translator_avalon_anti_slave_0_readdata;                                                      // uart_0:readdata -> uart_0_s1_translator:av_readdata
	wire         uart_0_s1_translator_avalon_anti_slave_0_begintransfer;                                                 // uart_0_s1_translator:av_begintransfer -> uart_0:begintransfer
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                               // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                 // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                     // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                      // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                  // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // SD_CMD_s1_translator:uav_waitrequest -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_CMD_s1_translator:uav_burstcount
	wire  [31:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_CMD_s1_translator:uav_writedata
	wire  [24:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_address -> SD_CMD_s1_translator:uav_address
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_write -> SD_CMD_s1_translator:uav_write
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SD_CMD_s1_translator:uav_lock
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_read -> SD_CMD_s1_translator:uav_read
	wire  [31:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // SD_CMD_s1_translator:uav_readdata -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // SD_CMD_s1_translator:uav_readdatavalid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_CMD_s1_translator:uav_debugaccess
	wire   [3:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_CMD_s1_translator:uav_byteenable
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // SD_DAT_s1_translator:uav_waitrequest -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_DAT_s1_translator:uav_burstcount
	wire  [31:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_DAT_s1_translator:uav_writedata
	wire  [24:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_address -> SD_DAT_s1_translator:uav_address
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_write -> SD_DAT_s1_translator:uav_write
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SD_DAT_s1_translator:uav_lock
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_read -> SD_DAT_s1_translator:uav_read
	wire  [31:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // SD_DAT_s1_translator:uav_readdata -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // SD_DAT_s1_translator:uav_readdatavalid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_DAT_s1_translator:uav_debugaccess
	wire   [3:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_DAT_s1_translator:uav_byteenable
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                  // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	wire  [24:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                   // nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // switch_pio_s1_translator:uav_waitrequest -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch_pio_s1_translator:uav_burstcount
	wire  [31:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch_pio_s1_translator:uav_writedata
	wire  [24:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch_pio_s1_translator:uav_address
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch_pio_s1_translator:uav_write
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch_pio_s1_translator:uav_lock
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch_pio_s1_translator:uav_read
	wire  [31:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // switch_pio_s1_translator:uav_readdata -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // switch_pio_s1_translator:uav_readdatavalid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch_pio_s1_translator:uav_debugaccess
	wire   [3:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch_pio_s1_translator:uav_byteenable
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	wire  [24:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	wire   [3:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // led_green_s1_translator:uav_waitrequest -> led_green_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led_green_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // led_green_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_green_s1_translator:uav_burstcount
	wire  [31:0] led_green_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // led_green_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_green_s1_translator:uav_writedata
	wire  [24:0] led_green_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // led_green_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_green_s1_translator:uav_address
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // led_green_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_green_s1_translator:uav_write
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // led_green_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_green_s1_translator:uav_lock
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // led_green_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_green_s1_translator:uav_read
	wire  [31:0] led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // led_green_s1_translator:uav_readdata -> led_green_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // led_green_s1_translator:uav_readdatavalid -> led_green_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // led_green_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_green_s1_translator:uav_debugaccess
	wire   [3:0] led_green_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // led_green_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_green_s1_translator:uav_byteenable
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // led_green_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // led_green_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // led_green_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // led_green_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_green_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // led_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led_red_s1_translator:uav_waitrequest -> led_red_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led_red_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led_red_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_red_s1_translator:uav_burstcount
	wire  [31:0] led_red_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led_red_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_red_s1_translator:uav_writedata
	wire  [24:0] led_red_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led_red_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_red_s1_translator:uav_address
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led_red_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_red_s1_translator:uav_write
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led_red_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_red_s1_translator:uav_lock
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led_red_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_red_s1_translator:uav_read
	wire  [31:0] led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led_red_s1_translator:uav_readdata -> led_red_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led_red_s1_translator:uav_readdatavalid -> led_red_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led_red_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_red_s1_translator:uav_debugaccess
	wire   [3:0] led_red_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led_red_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_red_s1_translator:uav_byteenable
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led_red_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led_red_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led_red_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led_red_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_red_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [24:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // cfi_flash_0_uas_translator:uav_waitrequest -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> cfi_flash_0_uas_translator:uav_burstcount
	wire   [7:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> cfi_flash_0_uas_translator:uav_writedata
	wire  [24:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address;                                   // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_address -> cfi_flash_0_uas_translator:uav_address
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write;                                     // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_write -> cfi_flash_0_uas_translator:uav_write
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                      // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_lock -> cfi_flash_0_uas_translator:uav_lock
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read;                                      // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_read -> cfi_flash_0_uas_translator:uav_read
	wire   [7:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // cfi_flash_0_uas_translator:uav_readdata -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // cfi_flash_0_uas_translator:uav_readdatavalid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cfi_flash_0_uas_translator:uav_debugaccess
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> cfi_flash_0_uas_translator:uav_byteenable
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [57:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                               // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [57:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // sram_16bit_512k_0_avalon_slave_0_translator:uav_waitrequest -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;               // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_16bit_512k_0_avalon_slave_0_translator:uav_burstcount
	wire  [15:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_16bit_512k_0_avalon_slave_0_translator:uav_writedata
	wire  [24:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                  // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> sram_16bit_512k_0_avalon_slave_0_translator:uav_address
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                    // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> sram_16bit_512k_0_avalon_slave_0_translator:uav_write
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                     // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> sram_16bit_512k_0_avalon_slave_0_translator:uav_lock
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                     // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> sram_16bit_512k_0_avalon_slave_0_translator:uav_read
	wire  [15:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                 // sram_16bit_512k_0_avalon_slave_0_translator:uav_readdata -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // sram_16bit_512k_0_avalon_slave_0_translator:uav_readdatavalid -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_16bit_512k_0_avalon_slave_0_translator:uav_debugaccess
	wire   [1:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;               // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_16bit_512k_0_avalon_slave_0_translator:uav_byteenable
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;             // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;              // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;             // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // sdram_0_s1_translator:uav_waitrequest -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_s1_translator:uav_burstcount
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_s1_translator:uav_writedata
	wire  [24:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_s1_translator:uav_address
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_s1_translator:uav_write
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_s1_translator:uav_lock
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_s1_translator:uav_read
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // sdram_0_s1_translator:uav_readdata -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // sdram_0_s1_translator:uav_readdatavalid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_s1_translator:uav_debugaccess
	wire   [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_s1_translator:uav_byteenable
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // epcs_controller_epcs_control_port_translator:uav_waitrequest -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;              // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> epcs_controller_epcs_control_port_translator:uav_burstcount
	wire  [31:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;               // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> epcs_controller_epcs_control_port_translator:uav_writedata
	wire  [24:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address;                 // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_address -> epcs_controller_epcs_control_port_translator:uav_address
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write;                   // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_write -> epcs_controller_epcs_control_port_translator:uav_write
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                    // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> epcs_controller_epcs_control_port_translator:uav_lock
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read;                    // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_read -> epcs_controller_epcs_control_port_translator:uav_read
	wire  [31:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                // epcs_controller_epcs_control_port_translator:uav_readdata -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // epcs_controller_epcs_control_port_translator:uav_readdatavalid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> epcs_controller_epcs_control_port_translator:uav_debugaccess
	wire   [3:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;              // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> epcs_controller_epcs_control_port_translator:uav_byteenable
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;            // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;             // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;            // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // uart_0_s1_translator:uav_waitrequest -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_0_s1_translator:uav_burstcount
	wire  [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_0_s1_translator:uav_writedata
	wire  [24:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_0_s1_translator:uav_address
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_0_s1_translator:uav_write
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_0_s1_translator:uav_lock
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_0_s1_translator:uav_read
	wire  [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // uart_0_s1_translator:uav_readdata -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // uart_0_s1_translator:uav_readdatavalid -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_0_s1_translator:uav_debugaccess
	wire   [3:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_0_s1_translator:uav_byteenable
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                       // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount;                        // nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata;                         // nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [24:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address;                           // nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock;                              // nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write;                             // nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read;                              // nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata;                          // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                       // nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable;                        // nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                     // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // SD_CLK_s1_translator:uav_waitrequest -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_CLK_s1_translator:uav_burstcount
	wire  [31:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_CLK_s1_translator:uav_writedata
	wire  [24:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_address -> SD_CLK_s1_translator:uav_address
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_write -> SD_CLK_s1_translator:uav_write
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SD_CLK_s1_translator:uav_lock
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_read -> SD_CLK_s1_translator:uav_read
	wire  [31:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // SD_CLK_s1_translator:uav_readdata -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // SD_CLK_s1_translator:uav_readdatavalid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_CLK_s1_translator:uav_debugaccess
	wire   [3:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_CLK_s1_translator:uav_byteenable
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // button_pio_s1_translator:uav_waitrequest -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_pio_s1_translator:uav_burstcount
	wire  [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_pio_s1_translator:uav_writedata
	wire  [24:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_pio_s1_translator:uav_address
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_pio_s1_translator:uav_write
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_pio_s1_translator:uav_lock
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_pio_s1_translator:uav_read
	wire  [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // button_pio_s1_translator:uav_readdata -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // button_pio_s1_translator:uav_readdatavalid -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_pio_s1_translator:uav_debugaccess
	wire   [3:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_pio_s1_translator:uav_byteenable
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // SEG7_Display_avalon_slave_translator:uav_waitrequest -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> SEG7_Display_avalon_slave_translator:uav_burstcount
	wire  [31:0] seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> SEG7_Display_avalon_slave_translator:uav_writedata
	wire  [24:0] seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> SEG7_Display_avalon_slave_translator:uav_address
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> SEG7_Display_avalon_slave_translator:uav_write
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> SEG7_Display_avalon_slave_translator:uav_lock
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> SEG7_Display_avalon_slave_translator:uav_read
	wire  [31:0] seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // SEG7_Display_avalon_slave_translator:uav_readdata -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // SEG7_Display_avalon_slave_translator:uav_readdatavalid -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SEG7_Display_avalon_slave_translator:uav_debugaccess
	wire   [3:0] seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> SEG7_Display_avalon_slave_translator:uav_byteenable
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest;                              // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount;                               // nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata;                                // nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [24:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_address;                                  // nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock;                                     // nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_write;                                    // nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_read;                                     // nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata;                                 // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess;                              // nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable;                               // nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid;                            // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [24:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                    // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // Audio_0_avalon_slave_0_translator:uav_waitrequest -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Audio_0_avalon_slave_0_translator:uav_burstcount
	wire  [31:0] audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                          // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Audio_0_avalon_slave_0_translator:uav_writedata
	wire  [24:0] audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                            // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Audio_0_avalon_slave_0_translator:uav_address
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                              // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Audio_0_avalon_slave_0_translator:uav_write
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                               // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Audio_0_avalon_slave_0_translator:uav_lock
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                               // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Audio_0_avalon_slave_0_translator:uav_read
	wire  [31:0] audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                           // Audio_0_avalon_slave_0_translator:uav_readdata -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // Audio_0_avalon_slave_0_translator:uav_readdatavalid -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Audio_0_avalon_slave_0_translator:uav_debugaccess
	wire   [3:0] audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Audio_0_avalon_slave_0_translator:uav_byteenable
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [84:0] audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                        // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [84:0] audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;              // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                    // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;            // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [83:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                     // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                    // addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                     // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                           // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                   // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [83:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                            // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                           // addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [83:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                    // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [65:0] sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                     // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_001:sink_ready -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                   // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [83:0] epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data;                    // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_002:sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                     // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [56:0] cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data;                                      // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_003:sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [65:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_004:sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                              // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [83:0] audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                               // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_005:sink_ready -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [83:0] seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_006:sink_ready -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // led_green_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // led_green_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // led_green_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [83:0] led_green_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // led_green_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         led_green_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_007:sink_ready -> led_green_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led_red_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led_red_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led_red_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [83:0] led_red_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led_red_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         led_red_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_008:sink_ready -> led_red_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [83:0] sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_009:sink_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [83:0] sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_010:sink_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [83:0] sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_011:sink_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [83:0] switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_012:sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [83:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_013:sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [83:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire         timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_014:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [83:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_015:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [83:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire         uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_016:sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [83:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_017:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                            // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                                  // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                          // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [83:0] addr_router_src_data;                                                                                   // addr_router:src_data -> limiter:cmd_sink_data
	wire  [17:0] addr_router_src_channel;                                                                                // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                                  // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                            // limiter:rsp_src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                                  // limiter:rsp_src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                          // limiter:rsp_src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [83:0] limiter_rsp_src_data;                                                                                   // limiter:rsp_src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [17:0] limiter_rsp_src_channel;                                                                                // limiter:rsp_src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                        // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                              // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                      // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [83:0] addr_router_001_src_data;                                                                               // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire  [17:0] addr_router_001_src_channel;                                                                            // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                              // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                        // limiter_001:rsp_src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                              // limiter_001:rsp_src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                      // limiter_001:rsp_src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [83:0] limiter_001_rsp_src_data;                                                                               // limiter_001:rsp_src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [17:0] limiter_001_rsp_src_channel;                                                                            // limiter_001:rsp_src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                              // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         burst_adapter_source0_endofpacket;                                                                      // burst_adapter:source0_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                            // burst_adapter:source0_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                                    // burst_adapter:source0_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [56:0] burst_adapter_source0_data;                                                                             // burst_adapter:source0_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                            // cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire  [17:0] burst_adapter_source0_channel;                                                                          // burst_adapter:source0_channel -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_001_source0_endofpacket;                                                                  // burst_adapter_001:source0_endofpacket -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_001_source0_valid;                                                                        // burst_adapter_001:source0_valid -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_001_source0_startofpacket;                                                                // burst_adapter_001:source0_startofpacket -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_001_source0_data;                                                                         // burst_adapter_001:source0_data -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_001_source0_ready;                                                                        // sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire  [17:0] burst_adapter_001_source0_channel;                                                                      // burst_adapter_001:source0_channel -> sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_002_source0_endofpacket;                                                                  // burst_adapter_002:source0_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_002_source0_valid;                                                                        // burst_adapter_002:source0_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_002_source0_startofpacket;                                                                // burst_adapter_002:source0_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_002_source0_data;                                                                         // burst_adapter_002:source0_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_002_source0_ready;                                                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire  [17:0] burst_adapter_002_source0_channel;                                                                      // burst_adapter_002:source0_channel -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rst_controller_reset_out_reset;                                                                         // rst_controller:reset_out -> [Audio_0:iRST_N, Audio_0_avalon_slave_0_translator:reset, Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_CLK:reset_n, SD_CLK_s1_translator:reset, SD_CLK_s1_translator_avalon_universal_slave_0_agent:reset, SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_CMD:reset_n, SD_CMD_s1_translator:reset, SD_CMD_s1_translator_avalon_universal_slave_0_agent:reset, SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_DAT:reset_n, SD_DAT_s1_translator:reset, SD_DAT_s1_translator_avalon_universal_slave_0_agent:reset, SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SEG7_Display:iRST_N, SEG7_Display_avalon_slave_translator:reset, SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:reset, SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, button_pio:reset_n, button_pio_s1_translator:reset, button_pio_s1_translator_avalon_universal_slave_0_agent:reset, button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cfi_flash_0:reset_reset, cfi_flash_0_uas_translator:reset, cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:reset, cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, epcs_controller:reset_n, epcs_controller_epcs_control_port_translator:reset, epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:reset, epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_green:reset_n, led_green_s1_translator:reset, led_green_s1_translator_avalon_universal_slave_0_agent:reset, led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_red:reset_n, led_red_s1_translator:reset, led_red_s1_translator_avalon_universal_slave_0_agent:reset, led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2_qsys_0:reset_n, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram_0:reset_n, sdram_0_s1_translator:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sram_16bit_512k_0:iRST_N, sram_16bit_512k_0_avalon_slave_0_translator:reset, sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch_pio:reset_n, switch_pio_s1_translator:reset, switch_pio_s1_translator_avalon_universal_slave_0_agent:reset, switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_1:reset_n, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tri_state_bridge_0_bridge_0:reset, tri_state_bridge_0_pinSharer_0:reset_reset, uart_0:reset_n, uart_0_s1_translator:reset, uart_0_s1_translator_avalon_universal_slave_0_agent:reset, uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                                                             // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         cmd_xbar_demux_src0_endofpacket;                                                                        // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                              // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                      // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [83:0] cmd_xbar_demux_src0_data;                                                                               // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [17:0] cmd_xbar_demux_src0_channel;                                                                            // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                              // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                        // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                              // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                      // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [83:0] cmd_xbar_demux_src1_data;                                                                               // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [17:0] cmd_xbar_demux_src1_channel;                                                                            // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                              // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                        // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                              // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                      // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [83:0] cmd_xbar_demux_src2_data;                                                                               // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [17:0] cmd_xbar_demux_src2_channel;                                                                            // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                              // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_src3_endofpacket;                                                                        // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                              // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                      // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [83:0] cmd_xbar_demux_src3_data;                                                                               // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire  [17:0] cmd_xbar_demux_src3_channel;                                                                            // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire         cmd_xbar_demux_src3_ready;                                                                              // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire         cmd_xbar_demux_src4_endofpacket;                                                                        // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                              // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                                      // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [83:0] cmd_xbar_demux_src4_data;                                                                               // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire  [17:0] cmd_xbar_demux_src4_channel;                                                                            // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire         cmd_xbar_demux_src4_ready;                                                                              // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                    // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                          // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                                  // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src0_data;                                                                           // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [17:0] cmd_xbar_demux_001_src0_channel;                                                                        // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                          // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                    // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                          // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                                  // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src1_data;                                                                           // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [17:0] cmd_xbar_demux_001_src1_channel;                                                                        // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                          // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                    // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                          // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                                  // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src2_data;                                                                           // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire  [17:0] cmd_xbar_demux_001_src2_channel;                                                                        // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                          // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                    // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                          // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                                  // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src3_data;                                                                           // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire  [17:0] cmd_xbar_demux_001_src3_channel;                                                                        // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire         cmd_xbar_demux_001_src3_ready;                                                                          // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                    // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                          // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                                  // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src4_data;                                                                           // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire  [17:0] cmd_xbar_demux_001_src4_channel;                                                                        // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire         cmd_xbar_demux_001_src4_ready;                                                                          // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                    // cmd_xbar_demux_001:src5_endofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                          // cmd_xbar_demux_001:src5_valid -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                                  // cmd_xbar_demux_001:src5_startofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src5_data;                                                                           // cmd_xbar_demux_001:src5_data -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src5_channel;                                                                        // cmd_xbar_demux_001:src5_channel -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                    // cmd_xbar_demux_001:src6_endofpacket -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                          // cmd_xbar_demux_001:src6_valid -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                                  // cmd_xbar_demux_001:src6_startofpacket -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src6_data;                                                                           // cmd_xbar_demux_001:src6_data -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src6_channel;                                                                        // cmd_xbar_demux_001:src6_channel -> SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                    // cmd_xbar_demux_001:src7_endofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                          // cmd_xbar_demux_001:src7_valid -> led_green_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                                  // cmd_xbar_demux_001:src7_startofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src7_data;                                                                           // cmd_xbar_demux_001:src7_data -> led_green_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src7_channel;                                                                        // cmd_xbar_demux_001:src7_channel -> led_green_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                    // cmd_xbar_demux_001:src8_endofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                          // cmd_xbar_demux_001:src8_valid -> led_red_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                                  // cmd_xbar_demux_001:src8_startofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src8_data;                                                                           // cmd_xbar_demux_001:src8_data -> led_red_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src8_channel;                                                                        // cmd_xbar_demux_001:src8_channel -> led_red_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                                    // cmd_xbar_demux_001:src9_endofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                          // cmd_xbar_demux_001:src9_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                                  // cmd_xbar_demux_001:src9_startofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src9_data;                                                                           // cmd_xbar_demux_001:src9_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src9_channel;                                                                        // cmd_xbar_demux_001:src9_channel -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                                   // cmd_xbar_demux_001:src10_endofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                         // cmd_xbar_demux_001:src10_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                                 // cmd_xbar_demux_001:src10_startofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src10_data;                                                                          // cmd_xbar_demux_001:src10_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src10_channel;                                                                       // cmd_xbar_demux_001:src10_channel -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src11_endofpacket;                                                                   // cmd_xbar_demux_001:src11_endofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src11_valid;                                                                         // cmd_xbar_demux_001:src11_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src11_startofpacket;                                                                 // cmd_xbar_demux_001:src11_startofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src11_data;                                                                          // cmd_xbar_demux_001:src11_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src11_channel;                                                                       // cmd_xbar_demux_001:src11_channel -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src12_endofpacket;                                                                   // cmd_xbar_demux_001:src12_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src12_valid;                                                                         // cmd_xbar_demux_001:src12_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src12_startofpacket;                                                                 // cmd_xbar_demux_001:src12_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src12_data;                                                                          // cmd_xbar_demux_001:src12_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src12_channel;                                                                       // cmd_xbar_demux_001:src12_channel -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src13_endofpacket;                                                                   // cmd_xbar_demux_001:src13_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src13_valid;                                                                         // cmd_xbar_demux_001:src13_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src13_startofpacket;                                                                 // cmd_xbar_demux_001:src13_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src13_data;                                                                          // cmd_xbar_demux_001:src13_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src13_channel;                                                                       // cmd_xbar_demux_001:src13_channel -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src14_endofpacket;                                                                   // cmd_xbar_demux_001:src14_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src14_valid;                                                                         // cmd_xbar_demux_001:src14_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src14_startofpacket;                                                                 // cmd_xbar_demux_001:src14_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src14_data;                                                                          // cmd_xbar_demux_001:src14_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src14_channel;                                                                       // cmd_xbar_demux_001:src14_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src15_endofpacket;                                                                   // cmd_xbar_demux_001:src15_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src15_valid;                                                                         // cmd_xbar_demux_001:src15_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src15_startofpacket;                                                                 // cmd_xbar_demux_001:src15_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src15_data;                                                                          // cmd_xbar_demux_001:src15_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src15_channel;                                                                       // cmd_xbar_demux_001:src15_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src16_endofpacket;                                                                   // cmd_xbar_demux_001:src16_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src16_valid;                                                                         // cmd_xbar_demux_001:src16_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src16_startofpacket;                                                                 // cmd_xbar_demux_001:src16_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src16_data;                                                                          // cmd_xbar_demux_001:src16_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src16_channel;                                                                       // cmd_xbar_demux_001:src16_channel -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src17_endofpacket;                                                                   // cmd_xbar_demux_001:src17_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src17_valid;                                                                         // cmd_xbar_demux_001:src17_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src17_startofpacket;                                                                 // cmd_xbar_demux_001:src17_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_demux_001_src17_data;                                                                          // cmd_xbar_demux_001:src17_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_demux_001_src17_channel;                                                                       // cmd_xbar_demux_001:src17_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                        // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                              // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                      // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [83:0] rsp_xbar_demux_src0_data;                                                                               // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [17:0] rsp_xbar_demux_src0_channel;                                                                            // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                              // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                        // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                              // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                      // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [83:0] rsp_xbar_demux_src1_data;                                                                               // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [17:0] rsp_xbar_demux_src1_channel;                                                                            // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                              // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                    // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                          // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                                  // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [83:0] rsp_xbar_demux_001_src0_data;                                                                           // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [17:0] rsp_xbar_demux_001_src0_channel;                                                                        // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                          // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                    // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                          // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                                  // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [83:0] rsp_xbar_demux_001_src1_data;                                                                           // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [17:0] rsp_xbar_demux_001_src1_channel;                                                                        // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                          // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                    // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                          // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                                  // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [83:0] rsp_xbar_demux_002_src0_data;                                                                           // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [17:0] rsp_xbar_demux_002_src0_channel;                                                                        // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                          // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                    // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                          // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                                  // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [83:0] rsp_xbar_demux_002_src1_data;                                                                           // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [17:0] rsp_xbar_demux_002_src1_channel;                                                                        // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                          // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                    // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                          // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                                  // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [83:0] rsp_xbar_demux_003_src0_data;                                                                           // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire  [17:0] rsp_xbar_demux_003_src0_channel;                                                                        // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                          // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_003_src1_endofpacket;                                                                    // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src1_valid;                                                                          // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src1_startofpacket;                                                                  // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [83:0] rsp_xbar_demux_003_src1_data;                                                                           // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire  [17:0] rsp_xbar_demux_003_src1_channel;                                                                        // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src1_ready;                                                                          // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                    // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                          // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                                  // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [83:0] rsp_xbar_demux_004_src0_data;                                                                           // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire  [17:0] rsp_xbar_demux_004_src0_channel;                                                                        // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                          // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_004_src1_endofpacket;                                                                    // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src1_valid;                                                                          // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src1_startofpacket;                                                                  // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [83:0] rsp_xbar_demux_004_src1_data;                                                                           // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire  [17:0] rsp_xbar_demux_004_src1_channel;                                                                        // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src1_ready;                                                                          // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                    // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                          // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                                  // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [83:0] rsp_xbar_demux_005_src0_data;                                                                           // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire  [17:0] rsp_xbar_demux_005_src0_channel;                                                                        // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                          // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                    // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                          // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                                  // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [83:0] rsp_xbar_demux_006_src0_data;                                                                           // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire  [17:0] rsp_xbar_demux_006_src0_channel;                                                                        // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                          // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                    // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                          // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                                  // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [83:0] rsp_xbar_demux_007_src0_data;                                                                           // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [17:0] rsp_xbar_demux_007_src0_channel;                                                                        // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                          // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                    // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                          // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                                  // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [83:0] rsp_xbar_demux_008_src0_data;                                                                           // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire  [17:0] rsp_xbar_demux_008_src0_channel;                                                                        // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                          // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                    // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                          // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                                  // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [83:0] rsp_xbar_demux_009_src0_data;                                                                           // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire  [17:0] rsp_xbar_demux_009_src0_channel;                                                                        // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                          // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                                    // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                          // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                                  // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [83:0] rsp_xbar_demux_010_src0_data;                                                                           // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire  [17:0] rsp_xbar_demux_010_src0_channel;                                                                        // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                          // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                                    // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                          // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                                  // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [83:0] rsp_xbar_demux_011_src0_data;                                                                           // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire  [17:0] rsp_xbar_demux_011_src0_channel;                                                                        // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                          // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                                    // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                          // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                                  // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [83:0] rsp_xbar_demux_012_src0_data;                                                                           // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire  [17:0] rsp_xbar_demux_012_src0_channel;                                                                        // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                          // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                                    // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                          // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                                  // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [83:0] rsp_xbar_demux_013_src0_data;                                                                           // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire  [17:0] rsp_xbar_demux_013_src0_channel;                                                                        // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                                          // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire         rsp_xbar_demux_014_src0_endofpacket;                                                                    // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire         rsp_xbar_demux_014_src0_valid;                                                                          // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire         rsp_xbar_demux_014_src0_startofpacket;                                                                  // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [83:0] rsp_xbar_demux_014_src0_data;                                                                           // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire  [17:0] rsp_xbar_demux_014_src0_channel;                                                                        // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire         rsp_xbar_demux_014_src0_ready;                                                                          // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire         rsp_xbar_demux_015_src0_endofpacket;                                                                    // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire         rsp_xbar_demux_015_src0_valid;                                                                          // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire         rsp_xbar_demux_015_src0_startofpacket;                                                                  // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [83:0] rsp_xbar_demux_015_src0_data;                                                                           // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire  [17:0] rsp_xbar_demux_015_src0_channel;                                                                        // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire         rsp_xbar_demux_015_src0_ready;                                                                          // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire         rsp_xbar_demux_016_src0_endofpacket;                                                                    // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire         rsp_xbar_demux_016_src0_valid;                                                                          // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire         rsp_xbar_demux_016_src0_startofpacket;                                                                  // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [83:0] rsp_xbar_demux_016_src0_data;                                                                           // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire  [17:0] rsp_xbar_demux_016_src0_channel;                                                                        // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire         rsp_xbar_demux_016_src0_ready;                                                                          // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire         rsp_xbar_demux_017_src0_endofpacket;                                                                    // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire         rsp_xbar_demux_017_src0_valid;                                                                          // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire         rsp_xbar_demux_017_src0_startofpacket;                                                                  // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [83:0] rsp_xbar_demux_017_src0_data;                                                                           // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire  [17:0] rsp_xbar_demux_017_src0_channel;                                                                        // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire         rsp_xbar_demux_017_src0_ready;                                                                          // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                            // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                          // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [83:0] limiter_cmd_src_data;                                                                                   // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire  [17:0] limiter_cmd_src_channel;                                                                                // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                                  // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                           // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                                 // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                         // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [83:0] rsp_xbar_mux_src_data;                                                                                  // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire  [17:0] rsp_xbar_mux_src_channel;                                                                               // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                                 // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                        // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                      // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [83:0] limiter_001_cmd_src_data;                                                                               // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire  [17:0] limiter_001_cmd_src_channel;                                                                            // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                              // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                       // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                             // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                     // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [83:0] rsp_xbar_mux_001_src_data;                                                                              // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire  [17:0] rsp_xbar_mux_001_src_channel;                                                                           // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                             // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                           // cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                                 // cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                         // cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_mux_src_data;                                                                                  // cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_mux_src_channel;                                                                               // cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                              // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                    // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                            // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [83:0] id_router_src_data;                                                                                     // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [17:0] id_router_src_channel;                                                                                  // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                    // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                       // cmd_xbar_mux_002:src_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                             // cmd_xbar_mux_002:src_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                     // cmd_xbar_mux_002:src_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [83:0] cmd_xbar_mux_002_src_data;                                                                              // cmd_xbar_mux_002:src_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire  [17:0] cmd_xbar_mux_002_src_channel;                                                                           // cmd_xbar_mux_002:src_channel -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                             // epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                          // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                                // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                        // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [83:0] id_router_002_src_data;                                                                                 // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [17:0] id_router_002_src_channel;                                                                              // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                                // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                          // Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                          // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                                // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                        // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [83:0] id_router_005_src_data;                                                                                 // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [17:0] id_router_005_src_channel;                                                                              // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                                // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                          // SEG7_Display_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                          // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                                // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                        // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [83:0] id_router_006_src_data;                                                                                 // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [17:0] id_router_006_src_channel;                                                                              // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                                // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                          // led_green_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                                          // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                                // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                        // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [83:0] id_router_007_src_data;                                                                                 // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [17:0] id_router_007_src_channel;                                                                              // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                                // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                          // led_red_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                          // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                                // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                        // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [83:0] id_router_008_src_data;                                                                                 // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [17:0] id_router_008_src_channel;                                                                              // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                                // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_demux_001_src9_ready;                                                                          // SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire         id_router_009_src_endofpacket;                                                                          // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                                // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                        // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [83:0] id_router_009_src_data;                                                                                 // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [17:0] id_router_009_src_channel;                                                                              // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                                // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_demux_001_src10_ready;                                                                         // SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire         id_router_010_src_endofpacket;                                                                          // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                                // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                        // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [83:0] id_router_010_src_data;                                                                                 // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [17:0] id_router_010_src_channel;                                                                              // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                                // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_demux_001_src11_ready;                                                                         // SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire         id_router_011_src_endofpacket;                                                                          // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                                // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                        // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [83:0] id_router_011_src_data;                                                                                 // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [17:0] id_router_011_src_channel;                                                                              // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                                // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         cmd_xbar_demux_001_src12_ready;                                                                         // switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire         id_router_012_src_endofpacket;                                                                          // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                                // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                        // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [83:0] id_router_012_src_data;                                                                                 // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [17:0] id_router_012_src_channel;                                                                              // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                                // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_demux_001_src13_ready;                                                                         // button_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire         id_router_013_src_endofpacket;                                                                          // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                                // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                        // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [83:0] id_router_013_src_data;                                                                                 // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire  [17:0] id_router_013_src_channel;                                                                              // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                                // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire         cmd_xbar_demux_001_src14_ready;                                                                         // timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire         id_router_014_src_endofpacket;                                                                          // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire         id_router_014_src_valid;                                                                                // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire         id_router_014_src_startofpacket;                                                                        // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [83:0] id_router_014_src_data;                                                                                 // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire  [17:0] id_router_014_src_channel;                                                                              // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire         id_router_014_src_ready;                                                                                // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire         cmd_xbar_demux_001_src15_ready;                                                                         // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire         id_router_015_src_endofpacket;                                                                          // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire         id_router_015_src_valid;                                                                                // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire         id_router_015_src_startofpacket;                                                                        // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [83:0] id_router_015_src_data;                                                                                 // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire  [17:0] id_router_015_src_channel;                                                                              // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire         id_router_015_src_ready;                                                                                // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire         cmd_xbar_demux_001_src16_ready;                                                                         // uart_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire         id_router_016_src_endofpacket;                                                                          // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire         id_router_016_src_valid;                                                                                // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire         id_router_016_src_startofpacket;                                                                        // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [83:0] id_router_016_src_data;                                                                                 // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire  [17:0] id_router_016_src_channel;                                                                              // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire         id_router_016_src_ready;                                                                                // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire         cmd_xbar_demux_001_src17_ready;                                                                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire         id_router_017_src_endofpacket;                                                                          // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire         id_router_017_src_valid;                                                                                // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire         id_router_017_src_startofpacket;                                                                        // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [83:0] id_router_017_src_data;                                                                                 // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire  [17:0] id_router_017_src_channel;                                                                              // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire         id_router_017_src_ready;                                                                                // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                       // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                             // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                     // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [83:0] cmd_xbar_mux_001_src_data;                                                                              // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire  [17:0] cmd_xbar_mux_001_src_channel;                                                                           // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                             // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire         width_adapter_src_endofpacket;                                                                          // width_adapter:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                                // width_adapter:out_valid -> burst_adapter_001:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                        // width_adapter:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [65:0] width_adapter_src_data;                                                                                 // width_adapter:out_data -> burst_adapter_001:sink0_data
	wire         width_adapter_src_ready;                                                                                // burst_adapter_001:sink0_ready -> width_adapter:out_ready
	wire  [17:0] width_adapter_src_channel;                                                                              // width_adapter:out_channel -> burst_adapter_001:sink0_channel
	wire         id_router_001_src_endofpacket;                                                                          // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_001_src_valid;                                                                                // id_router_001:src_valid -> width_adapter_001:in_valid
	wire         id_router_001_src_startofpacket;                                                                        // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [65:0] id_router_001_src_data;                                                                                 // id_router_001:src_data -> width_adapter_001:in_data
	wire  [17:0] id_router_001_src_channel;                                                                              // id_router_001:src_channel -> width_adapter_001:in_channel
	wire         id_router_001_src_ready;                                                                                // width_adapter_001:in_ready -> id_router_001:src_ready
	wire         width_adapter_001_src_endofpacket;                                                                      // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                                            // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                                    // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [83:0] width_adapter_001_src_data;                                                                             // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire         width_adapter_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire  [17:0] width_adapter_001_src_channel;                                                                          // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire         cmd_xbar_mux_003_src_endofpacket;                                                                       // cmd_xbar_mux_003:src_endofpacket -> width_adapter_002:in_endofpacket
	wire         cmd_xbar_mux_003_src_valid;                                                                             // cmd_xbar_mux_003:src_valid -> width_adapter_002:in_valid
	wire         cmd_xbar_mux_003_src_startofpacket;                                                                     // cmd_xbar_mux_003:src_startofpacket -> width_adapter_002:in_startofpacket
	wire  [83:0] cmd_xbar_mux_003_src_data;                                                                              // cmd_xbar_mux_003:src_data -> width_adapter_002:in_data
	wire  [17:0] cmd_xbar_mux_003_src_channel;                                                                           // cmd_xbar_mux_003:src_channel -> width_adapter_002:in_channel
	wire         cmd_xbar_mux_003_src_ready;                                                                             // width_adapter_002:in_ready -> cmd_xbar_mux_003:src_ready
	wire         width_adapter_002_src_endofpacket;                                                                      // width_adapter_002:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_002_src_valid;                                                                            // width_adapter_002:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_002_src_startofpacket;                                                                    // width_adapter_002:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [56:0] width_adapter_002_src_data;                                                                             // width_adapter_002:out_data -> burst_adapter:sink0_data
	wire         width_adapter_002_src_ready;                                                                            // burst_adapter:sink0_ready -> width_adapter_002:out_ready
	wire  [17:0] width_adapter_002_src_channel;                                                                          // width_adapter_002:out_channel -> burst_adapter:sink0_channel
	wire         id_router_003_src_endofpacket;                                                                          // id_router_003:src_endofpacket -> width_adapter_003:in_endofpacket
	wire         id_router_003_src_valid;                                                                                // id_router_003:src_valid -> width_adapter_003:in_valid
	wire         id_router_003_src_startofpacket;                                                                        // id_router_003:src_startofpacket -> width_adapter_003:in_startofpacket
	wire  [56:0] id_router_003_src_data;                                                                                 // id_router_003:src_data -> width_adapter_003:in_data
	wire  [17:0] id_router_003_src_channel;                                                                              // id_router_003:src_channel -> width_adapter_003:in_channel
	wire         id_router_003_src_ready;                                                                                // width_adapter_003:in_ready -> id_router_003:src_ready
	wire         width_adapter_003_src_endofpacket;                                                                      // width_adapter_003:out_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         width_adapter_003_src_valid;                                                                            // width_adapter_003:out_valid -> rsp_xbar_demux_003:sink_valid
	wire         width_adapter_003_src_startofpacket;                                                                    // width_adapter_003:out_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [83:0] width_adapter_003_src_data;                                                                             // width_adapter_003:out_data -> rsp_xbar_demux_003:sink_data
	wire         width_adapter_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> width_adapter_003:out_ready
	wire  [17:0] width_adapter_003_src_channel;                                                                          // width_adapter_003:out_channel -> rsp_xbar_demux_003:sink_channel
	wire         cmd_xbar_mux_004_src_endofpacket;                                                                       // cmd_xbar_mux_004:src_endofpacket -> width_adapter_004:in_endofpacket
	wire         cmd_xbar_mux_004_src_valid;                                                                             // cmd_xbar_mux_004:src_valid -> width_adapter_004:in_valid
	wire         cmd_xbar_mux_004_src_startofpacket;                                                                     // cmd_xbar_mux_004:src_startofpacket -> width_adapter_004:in_startofpacket
	wire  [83:0] cmd_xbar_mux_004_src_data;                                                                              // cmd_xbar_mux_004:src_data -> width_adapter_004:in_data
	wire  [17:0] cmd_xbar_mux_004_src_channel;                                                                           // cmd_xbar_mux_004:src_channel -> width_adapter_004:in_channel
	wire         cmd_xbar_mux_004_src_ready;                                                                             // width_adapter_004:in_ready -> cmd_xbar_mux_004:src_ready
	wire         width_adapter_004_src_endofpacket;                                                                      // width_adapter_004:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire         width_adapter_004_src_valid;                                                                            // width_adapter_004:out_valid -> burst_adapter_002:sink0_valid
	wire         width_adapter_004_src_startofpacket;                                                                    // width_adapter_004:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire  [65:0] width_adapter_004_src_data;                                                                             // width_adapter_004:out_data -> burst_adapter_002:sink0_data
	wire         width_adapter_004_src_ready;                                                                            // burst_adapter_002:sink0_ready -> width_adapter_004:out_ready
	wire  [17:0] width_adapter_004_src_channel;                                                                          // width_adapter_004:out_channel -> burst_adapter_002:sink0_channel
	wire         id_router_004_src_endofpacket;                                                                          // id_router_004:src_endofpacket -> width_adapter_005:in_endofpacket
	wire         id_router_004_src_valid;                                                                                // id_router_004:src_valid -> width_adapter_005:in_valid
	wire         id_router_004_src_startofpacket;                                                                        // id_router_004:src_startofpacket -> width_adapter_005:in_startofpacket
	wire  [65:0] id_router_004_src_data;                                                                                 // id_router_004:src_data -> width_adapter_005:in_data
	wire  [17:0] id_router_004_src_channel;                                                                              // id_router_004:src_channel -> width_adapter_005:in_channel
	wire         id_router_004_src_ready;                                                                                // width_adapter_005:in_ready -> id_router_004:src_ready
	wire         width_adapter_005_src_endofpacket;                                                                      // width_adapter_005:out_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         width_adapter_005_src_valid;                                                                            // width_adapter_005:out_valid -> rsp_xbar_demux_004:sink_valid
	wire         width_adapter_005_src_startofpacket;                                                                    // width_adapter_005:out_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [83:0] width_adapter_005_src_data;                                                                             // width_adapter_005:out_data -> rsp_xbar_demux_004:sink_data
	wire         width_adapter_005_src_ready;                                                                            // rsp_xbar_demux_004:sink_ready -> width_adapter_005:out_ready
	wire  [17:0] width_adapter_005_src_channel;                                                                          // width_adapter_005:out_channel -> rsp_xbar_demux_004:sink_channel
	wire  [17:0] limiter_cmd_valid_data;                                                                                 // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire  [17:0] limiter_001_cmd_valid_data;                                                                             // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                               // epcs_controller:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                               // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                               // uart_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                                               // timer_0:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                                               // button_pio:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                                               // timer_1:irq -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                                                                 // irq_mapper:sender_irq -> nios2_qsys_0:d_irq

	system_0_sdram_0 sdram_0 (
		.clk            (clk_clk_in_clk),                                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                         // reset.reset_n
		.az_addr        (sdram_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_0_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_0_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_0_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_0_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_0_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_0_wire_dq),                                         //      .export
		.zs_dqm         (sdram_0_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_0_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_0_wire_we_n)                                        //      .export
	);

	system_0_epcs_controller epcs_controller (
		.clk           (clk_clk_in_clk),                                                              //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                             //             reset.reset_n
		.address       (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address),    // epcs_control_port.address
		.chipselect    (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect), //                  .chipselect
		.dataavailable (),                                                                            //                  .dataavailable
		.endofpacket   (),                                                                            //                  .endofpacket
		.read_n        (~epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read),      //                  .read_n
		.readdata      (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata),   //                  .readdata
		.readyfordata  (),                                                                            //                  .readyfordata
		.write_n       (~epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write),     //                  .write_n
		.writedata     (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver0_irq)                                                     //               irq.irq
	);

	system_0_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk_in_clk),                                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.dataavailable  (),                                                                         //                  .dataavailable
		.readyfordata   (),                                                                         //                  .readyfordata
		.av_irq         (irq_mapper_receiver1_irq)                                                  //               irq.irq
	);

	system_0_uart_0 uart_0 (
		.clk           (clk_clk_in_clk),                                         //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address       (uart_0_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart_0_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart_0_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart_0_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart_0_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart_0_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart_0_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                       //                    .dataavailable
		.readyfordata  (),                                                       //                    .readyfordata
		.rxd           (uart_0_external_connection_rxd),                         // external_connection.export
		.txd           (uart_0_external_connection_txd),                         //                    .export
		.irq           (irq_mapper_receiver2_irq)                                //                 irq.irq
	);

	system_0_timer_0 timer_0 (
		.clk        (clk_clk_in_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                              //   irq.irq
	);

	system_0_timer_0 timer_1 (
		.clk        (clk_clk_in_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                              //   irq.irq
	);

	system_0_led_red led_red (
		.clk        (clk_clk_in_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (led_red_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_red_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_red_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_red_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_red_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_red_external_connection_export)                    // external_connection.export
	);

	system_0_led_green led_green (
		.clk        (clk_clk_in_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (led_green_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_green_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_green_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_green_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_green_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_green_external_connection_export)                    // external_connection.export
	);

	system_0_button_pio button_pio (
		.clk        (clk_clk_in_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (button_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~button_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (button_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (button_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (button_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (button_pio_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                                 //                 irq.irq
	);

	system_0_switch_pio switch_pio (
		.clk      (clk_clk_in_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address  (switch_pio_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (switch_pio_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (switch_pio_external_connection_export)                  // external_connection.export
	);

	system_0_SD_DAT sd_dat (
		.clk        (clk_clk_in_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (sd_dat_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sd_dat_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sd_dat_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sd_dat_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sd_dat_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (sd_dat_external_connection_export)                    // external_connection.export
	);

	system_0_SD_DAT sd_cmd (
		.clk        (clk_clk_in_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (sd_cmd_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sd_cmd_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sd_cmd_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sd_cmd_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sd_cmd_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (sd_cmd_external_connection_export)                    // external_connection.export
	);

	system_0_SD_CLK sd_clk (
		.clk        (clk_clk_in_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (sd_clk_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sd_clk_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sd_clk_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sd_clk_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sd_clk_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (sd_clk_external_connection_export)                    // external_connection.export
	);

	system_0_tri_state_bridge_0_bridge_0 tri_state_bridge_0_bridge_0 (
		.clk                               (clk_clk_in_clk),                                                     //   clk.clk
		.reset                             (rst_controller_reset_out_reset),                                     // reset.reset
		.request                           (tri_state_bridge_0_pinsharer_0_tcm_request),                         //   tcs.request
		.grant                             (tri_state_bridge_0_pinsharer_0_tcm_grant),                           //      .grant
		.tcs_tri_state_bridge_0_data       (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out),     //      .tri_state_bridge_0_data_out
		.tcs_tri_state_bridge_0_data_outen (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen),   //      .tri_state_bridge_0_data_outen
		.tcs_tri_state_bridge_0_data_in    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in),      //      .tri_state_bridge_0_data_in
		.tcs_tri_state_bridge_0_readn      (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out),    //      .tri_state_bridge_0_readn_out
		.tcs_write_n_to_the_cfi_flash_0    (tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out),  //      .write_n_to_the_cfi_flash_0_out
		.tcs_tri_state_bridge_0_address    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out),  //      .tri_state_bridge_0_address_out
		.tcs_select_n_to_the_cfi_flash_0   (tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out), //      .select_n_to_the_cfi_flash_0_out
		.tri_state_bridge_0_data           (tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_data),            //   out.tri_state_bridge_0_data
		.tri_state_bridge_0_readn          (tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_readn),           //      .tri_state_bridge_0_readn
		.write_n_to_the_cfi_flash_0        (tri_state_bridge_0_bridge_0_out_write_n_to_the_cfi_flash_0),         //      .write_n_to_the_cfi_flash_0
		.tri_state_bridge_0_address        (tri_state_bridge_0_bridge_0_out_tri_state_bridge_0_address),         //      .tri_state_bridge_0_address
		.select_n_to_the_cfi_flash_0       (tri_state_bridge_0_bridge_0_out_select_n_to_the_cfi_flash_0)         //      .select_n_to_the_cfi_flash_0
	);

	system_0_tri_state_bridge_0_pinSharer_0 tri_state_bridge_0_pinsharer_0 (
		.clk_clk                       (clk_clk_in_clk),                                                     //   clk.clk
		.reset_reset                   (rst_controller_reset_out_reset),                                     // reset.reset
		.request                       (tri_state_bridge_0_pinsharer_0_tcm_request),                         //   tcm.request
		.grant                         (tri_state_bridge_0_pinsharer_0_tcm_grant),                           //      .grant
		.tri_state_bridge_0_address    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out),  //      .tri_state_bridge_0_address_out
		.tri_state_bridge_0_readn      (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out),    //      .tri_state_bridge_0_readn_out
		.write_n_to_the_cfi_flash_0    (tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out),  //      .write_n_to_the_cfi_flash_0_out
		.tri_state_bridge_0_data       (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out),     //      .tri_state_bridge_0_data_out
		.tri_state_bridge_0_data_in    (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in),      //      .tri_state_bridge_0_data_in
		.tri_state_bridge_0_data_outen (tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen),   //      .tri_state_bridge_0_data_outen
		.select_n_to_the_cfi_flash_0   (tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out), //      .select_n_to_the_cfi_flash_0_out
		.tcs0_request                  (cfi_flash_0_tcm_request),                                            //  tcs0.request
		.tcs0_grant                    (cfi_flash_0_tcm_grant),                                              //      .grant
		.tcs0_address_out              (cfi_flash_0_tcm_address_out),                                        //      .address_out
		.tcs0_read_n_out               (cfi_flash_0_tcm_read_n_out),                                         //      .read_n_out
		.tcs0_write_n_out              (cfi_flash_0_tcm_write_n_out),                                        //      .write_n_out
		.tcs0_data_out                 (cfi_flash_0_tcm_data_out),                                           //      .data_out
		.tcs0_data_in                  (cfi_flash_0_tcm_data_in),                                            //      .data_in
		.tcs0_data_outen               (cfi_flash_0_tcm_data_outen),                                         //      .data_outen
		.tcs0_chipselect_n_out         (cfi_flash_0_tcm_chipselect_n_out)                                    //      .chipselect_n_out
	);

	system_0_cfi_flash_0 #(
		.TCM_ADDRESS_W                  (22),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (40),
		.TCM_DATA_HOLD                  (40),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) cfi_flash_0 (
		.clk_clk              (clk_clk_in_clk),                                               //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                               // reset.reset
		.uas_address          (cfi_flash_0_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (cfi_flash_0_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (cfi_flash_0_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (cfi_flash_0_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (cfi_flash_0_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (cfi_flash_0_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (cfi_flash_0_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (cfi_flash_0_tcm_request),                                      //      .request
		.tcm_grant            (cfi_flash_0_tcm_grant),                                        //      .grant
		.tcm_address_out      (cfi_flash_0_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (cfi_flash_0_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (cfi_flash_0_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (cfi_flash_0_tcm_data_in)                                       //      .data_in
	);

	SEG7_LUT_8 seg7_display (
		.iCLK   (clk_clk_in_clk),                                                     //          clk.clk
		.iWR    (seg7_display_avalon_slave_translator_avalon_anti_slave_0_write),     // avalon_slave.write
		.iDIG   (seg7_display_avalon_slave_translator_avalon_anti_slave_0_writedata), //             .writedata
		.oSEG0  (seg7_display_conduit_end_oSEG0),                                     //  conduit_end.export
		.oSEG1  (seg7_display_conduit_end_oSEG1),                                     //             .export
		.oSEG2  (seg7_display_conduit_end_oSEG2),                                     //             .export
		.oSEG3  (seg7_display_conduit_end_oSEG3),                                     //             .export
		.oSEG4  (seg7_display_conduit_end_oSEG4),                                     //             .export
		.oSEG5  (seg7_display_conduit_end_oSEG5),                                     //             .export
		.oSEG6  (seg7_display_conduit_end_oSEG6),                                     //             .export
		.oSEG7  (seg7_display_conduit_end_oSEG7),                                     //             .export
		.iRST_N (~rst_controller_reset_out_reset)                                     //      reset_n.reset_n
	);

	AUDIO_DAC_FIFO #(
		.REF_CLK     (18432000),
		.SAMPLE_RATE (48000),
		.DATA_WIDTH  (16),
		.CHANNEL_NUM (2)
	) audio_0 (
		.iWR_CLK   (clk_clk_in_clk),                                                  //                   clk.clk
		.oAUD_DATA (audio_0_avalon_slave_0_export_oAUD_DATA),                         // avalon_slave_0_export.export
		.oAUD_LRCK (audio_0_avalon_slave_0_export_oAUD_LRCK),                         //                      .export
		.oAUD_BCK  (audio_0_avalon_slave_0_export_oAUD_BCK),                          //                      .export
		.oAUD_XCK  (audio_0_avalon_slave_0_export_oAUD_XCK),                          //                      .export
		.iCLK_18_4 (audio_0_avalon_slave_0_export_iCLK_18_4),                         //                      .export
		.iDATA     (audio_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata), //        avalon_slave_0.writedata
		.iWR       (audio_0_avalon_slave_0_translator_avalon_anti_slave_0_write),     //                      .write
		.oDATA     (audio_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.iRST_N    (~rst_controller_reset_out_reset)                                  //               reset_n.reset_n
	);

	SRAM_16Bit_512K sram_16bit_512k_0 (
		.iCLK      (clk_clk_in_clk),                                                              //                   clk.clk
		.SRAM_DQ   (sram_16bit_512k_0_avalon_slave_0_export_DQ),                                  // avalon_slave_0_export.export
		.SRAM_ADDR (sram_16bit_512k_0_avalon_slave_0_export_ADDR),                                //                      .export
		.SRAM_UB_N (sram_16bit_512k_0_avalon_slave_0_export_UB_N),                                //                      .export
		.SRAM_LB_N (sram_16bit_512k_0_avalon_slave_0_export_LB_N),                                //                      .export
		.SRAM_WE_N (sram_16bit_512k_0_avalon_slave_0_export_WE_N),                                //                      .export
		.SRAM_CE_N (sram_16bit_512k_0_avalon_slave_0_export_CE_N),                                //                      .export
		.SRAM_OE_N (sram_16bit_512k_0_avalon_slave_0_export_OE_N),                                //                      .export
		.iDATA     (sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //        avalon_slave_0.writedata
		.oDATA     (sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //                      .readdata
		.iADDR     (sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_address),     //                      .address
		.iWE_N     (~sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //                      .write_n
		.iOE_N     (~sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       //                      .read_n
		.iCE_N     (~sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //                      .chipselect_n
		.iBE_N     (~sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //                      .byteenable_n
		.iRST_N    (~rst_controller_reset_out_reset)                                              //               reset_n.reset_n
	);

	system_0_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk_in_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                             //                   reset_n.reset_n
		.d_address                             (nios2_qsys_0_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (nios2_qsys_0_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                             // custom_instruction_master.readra
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_instruction_master_translator (
		.clk                   (clk_clk_in_clk),                                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_qsys_0_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_0_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_qsys_0_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                                               //               (terminated)
		.av_write              (1'b0),                                                                               //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock               (1'b0),                                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                                               //               (terminated)
		.uav_clken             (),                                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_data_master_translator (
		.clk                   (clk_clk_in_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_qsys_0_data_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_qsys_0_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (nios2_qsys_0_data_master_write),                                              //                          .write
		.av_writedata          (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_0_jtag_debug_module_translator (
		.clk                   (clk_clk_in_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                                          //              (terminated)
		.av_burstcount         (),                                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                                          //              (terminated)
		.av_lock               (),                                                                                          //              (terminated)
		.av_clken              (),                                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (2),
		.AV_WRITE_WAIT_CYCLES           (2),
		.AV_SETUP_WAIT_CYCLES           (2),
		.AV_DATA_HOLD_CYCLES            (2)
	) sram_16bit_512k_0_avalon_slave_0_translator (
		.clk                   (clk_clk_in_clk),                                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                              //                    reset.reset
		.uav_address           (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (sram_16bit_512k_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                                            //              (terminated)
		.av_burstcount         (),                                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                                            //              (terminated)
		.av_lock               (),                                                                                            //              (terminated)
		.av_clken              (),                                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                                        //              (terminated)
		.av_debugaccess        (),                                                                                            //              (terminated)
		.av_outputenable       ()                                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) epcs_controller_epcs_control_port_translator (
		.clk                   (clk_clk_in_clk),                                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                               //                    reset.reset
		.uav_address           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                             //              (terminated)
		.av_byteenable         (),                                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_lock               (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_debugaccess        (),                                                                                             //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cfi_flash_0_uas_translator (
		.clk                   (clk_clk_in_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                             //                    reset.reset
		.uav_address           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cfi_flash_0_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cfi_flash_0_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (cfi_flash_0_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (cfi_flash_0_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_chipselect         (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_0_s1_translator (
		.clk                   (clk_clk_in_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_0_avalon_slave_0_translator (
		.clk                   (clk_clk_in_clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (audio_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_readdata           (audio_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (audio_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_address            (),                                                                                  //              (terminated)
		.av_read               (),                                                                                  //              (terminated)
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_chipselect         (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seg7_display_avalon_slave_translator (
		.clk                   (clk_clk_in_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (seg7_display_avalon_slave_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (seg7_display_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_address            (),                                                                                     //              (terminated)
		.av_read               (),                                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                                 //              (terminated)
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                     //              (terminated)
		.av_byteenable         (),                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_chipselect         (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_green_s1_translator (
		.clk                   (clk_clk_in_clk),                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (led_green_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (led_green_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (led_green_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (led_green_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (led_green_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (led_green_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (led_green_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (led_green_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (led_green_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (led_green_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (led_green_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (led_green_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (led_green_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (led_green_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_red_s1_translator (
		.clk                   (clk_clk_in_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (led_red_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (led_red_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (led_red_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (led_red_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (led_red_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (led_red_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (led_red_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (led_red_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (led_red_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (led_red_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (led_red_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (led_red_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (led_red_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (led_red_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_clk_s1_translator (
		.clk                   (clk_clk_in_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_clk_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_clk_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sd_clk_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_clk_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sd_clk_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_cmd_s1_translator (
		.clk                   (clk_clk_in_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_cmd_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_cmd_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sd_cmd_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_cmd_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sd_cmd_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_dat_s1_translator (
		.clk                   (clk_clk_in_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sd_dat_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sd_dat_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sd_dat_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sd_dat_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sd_dat_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch_pio_s1_translator (
		.clk                   (clk_clk_in_clk),                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (switch_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (switch_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                         //              (terminated)
		.av_read               (),                                                                         //              (terminated)
		.av_writedata          (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button_pio_s1_translator (
		.clk                   (clk_clk_in_clk),                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (button_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (button_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (button_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (button_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (button_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_1_s1_translator (
		.clk                   (clk_clk_in_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                   (clk_clk_in_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_0_s1_translator (
		.clk                   (clk_clk_in_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (uart_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (uart_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (uart_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (uart_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (uart_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (uart_0_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect         (uart_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (clk_clk_in_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_cmd_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                               //                .channel
		.rf_sink_ready           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_dat_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                               //                .channel
		.rf_sink_ready           (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                            //                .channel
		.rf_sink_ready           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) switch_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                   //                .channel
		.rf_sink_ready           (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                                //                .channel
		.rf_sink_ready           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) led_green_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (led_green_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_green_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_green_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_green_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_green_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_green_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_green_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_green_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_green_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_green_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_green_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_green_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_green_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_green_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                   //                .channel
		.rf_sink_ready           (led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) led_red_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (led_red_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_red_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_red_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_red_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_red_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_red_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_red_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_red_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_red_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_red_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_red_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_red_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_red_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_red_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                 //                .channel
		.rf_sink_ready           (led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                                //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (45),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_POSTED          (35),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.PKT_TRANS_LOCK            (38),
		.PKT_SRC_ID_H              (50),
		.PKT_SRC_ID_L              (46),
		.PKT_DEST_ID_H             (55),
		.PKT_DEST_ID_L             (51),
		.PKT_BURSTWRAP_H           (44),
		.PKT_BURSTWRAP_L           (42),
		.PKT_BYTE_CNT_H            (41),
		.PKT_BYTE_CNT_L            (39),
		.PKT_PROTECTION_H          (56),
		.PKT_PROTECTION_L          (56),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (57),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cfi_flash_0_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                          //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                          //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                           //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                    //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                        //                .channel
		.rf_sink_ready           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (58),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (54),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (59),
		.PKT_SRC_ID_L              (55),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (60),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                                       //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                                       //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                        //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (54),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (59),
		.PKT_SRC_ID_L              (55),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (60),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                 //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                 //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                  //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                           //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                               //                .channel
		.rf_sink_ready           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                         //       clk_reset.reset
		.m0_address              (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                           //                .channel
		.rf_sink_ready           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                         // clk_reset.reset
		.in_data           (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) uart_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                               //                .channel
		.rf_sink_ready           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.PKT_BEGIN_BURST           (72),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (18),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3)
	) nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk_in_clk),                                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                       //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                        //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                                     //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                               //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                                 //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                        //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sd_clk_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                //                .channel
		.rf_sink_ready           (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) button_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                   //                .channel
		.rf_sink_ready           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                                //                .channel
		.rf_sink_ready           (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.PKT_BEGIN_BURST           (72),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (18),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7)
	) nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk_in_clk),                                                                       //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                                                   //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (77),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (83),
		.ST_CHANNEL_W              (18),
		.ST_DATA_W                 (84),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk_in_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                             //                .channel
		.rf_sink_ready           (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (85),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk_in_clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	system_0_addr_router addr_router (
		.sink_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                                       //          .valid
		.src_data           (addr_router_src_data),                                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                  //          .endofpacket
	);

	system_0_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	system_0_id_router id_router (
		.sink_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_src_valid),                                                                       //          .valid
		.src_data           (id_router_src_data),                                                                        //          .data
		.src_channel        (id_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                  //          .endofpacket
	);

	system_0_id_router_001 id_router_001 (
		.sink_ready         (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_16bit_512k_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_001_src_valid),                                                                     //          .valid
		.src_data           (id_router_001_src_data),                                                                      //          .data
		.src_channel        (id_router_001_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                                //          .endofpacket
	);

	system_0_id_router id_router_002 (
		.sink_ready         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                      //          .valid
		.src_data           (id_router_002_src_data),                                                                       //          .data
		.src_channel        (id_router_002_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                                 //          .endofpacket
	);

	system_0_id_router_003 id_router_003 (
		.sink_ready         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                    //       src.ready
		.src_valid          (id_router_003_src_valid),                                                    //          .valid
		.src_data           (id_router_003_src_data),                                                     //          .data
		.src_channel        (id_router_003_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                               //          .endofpacket
	);

	system_0_id_router_001 id_router_004 (
		.sink_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                               //       src.ready
		.src_valid          (id_router_004_src_valid),                                               //          .valid
		.src_data           (id_router_004_src_data),                                                //          .data
		.src_channel        (id_router_004_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_005 id_router_005 (
		.sink_ready         (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                           //       src.ready
		.src_valid          (id_router_005_src_valid),                                                           //          .valid
		.src_data           (id_router_005_src_data),                                                            //          .data
		.src_channel        (id_router_005_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                      //          .endofpacket
	);

	system_0_id_router_005 id_router_006 (
		.sink_ready         (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seg7_display_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                              //       src.ready
		.src_valid          (id_router_006_src_valid),                                                              //          .valid
		.src_data           (id_router_006_src_data),                                                               //          .data
		.src_channel        (id_router_006_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                         //          .endofpacket
	);

	system_0_id_router_005 id_router_007 (
		.sink_ready         (led_green_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_green_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_green_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_green_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_green_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                 //       src.ready
		.src_valid          (id_router_007_src_valid),                                                 //          .valid
		.src_data           (id_router_007_src_data),                                                  //          .data
		.src_channel        (id_router_007_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                            //          .endofpacket
	);

	system_0_id_router_005 id_router_008 (
		.sink_ready         (led_red_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_red_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_red_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_red_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_red_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                               //       src.ready
		.src_valid          (id_router_008_src_valid),                                               //          .valid
		.src_data           (id_router_008_src_data),                                                //          .data
		.src_channel        (id_router_008_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_005 id_router_009 (
		.sink_ready         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                              //       src.ready
		.src_valid          (id_router_009_src_valid),                                              //          .valid
		.src_data           (id_router_009_src_data),                                               //          .data
		.src_channel        (id_router_009_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                         //          .endofpacket
	);

	system_0_id_router_005 id_router_010 (
		.sink_ready         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                              //       src.ready
		.src_valid          (id_router_010_src_valid),                                              //          .valid
		.src_data           (id_router_010_src_data),                                               //          .data
		.src_channel        (id_router_010_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                         //          .endofpacket
	);

	system_0_id_router_005 id_router_011 (
		.sink_ready         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                              //       src.ready
		.src_valid          (id_router_011_src_valid),                                              //          .valid
		.src_data           (id_router_011_src_data),                                               //          .data
		.src_channel        (id_router_011_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                         //          .endofpacket
	);

	system_0_id_router_005 id_router_012 (
		.sink_ready         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                  //       src.ready
		.src_valid          (id_router_012_src_valid),                                                  //          .valid
		.src_data           (id_router_012_src_data),                                                   //          .data
		.src_channel        (id_router_012_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                             //          .endofpacket
	);

	system_0_id_router_005 id_router_013 (
		.sink_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                  //       src.ready
		.src_valid          (id_router_013_src_valid),                                                  //          .valid
		.src_data           (id_router_013_src_data),                                                   //          .data
		.src_channel        (id_router_013_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                             //          .endofpacket
	);

	system_0_id_router_005 id_router_014 (
		.sink_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                               //       src.ready
		.src_valid          (id_router_014_src_valid),                                               //          .valid
		.src_data           (id_router_014_src_data),                                                //          .data
		.src_channel        (id_router_014_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_005 id_router_015 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                               //       src.ready
		.src_valid          (id_router_015_src_valid),                                               //          .valid
		.src_data           (id_router_015_src_data),                                                //          .data
		.src_channel        (id_router_015_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                          //          .endofpacket
	);

	system_0_id_router_005 id_router_016 (
		.sink_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                              //       src.ready
		.src_valid          (id_router_016_src_valid),                                              //          .valid
		.src_data           (id_router_016_src_data),                                               //          .data
		.src_channel        (id_router_016_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                         //          .endofpacket
	);

	system_0_id_router_005 id_router_017 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk_in_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_017_src_valid),                                                                  //          .valid
		.src_data           (id_router_017_src_data),                                                                   //          .data
		.src_channel        (id_router_017_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                             //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_TRANS_POSTED          (62),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (18),
		.VALID_WIDTH               (18),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk_in_clk),                 //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (78),
		.PKT_TRANS_POSTED          (62),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (84),
		.ST_CHANNEL_W              (18),
		.VALID_WIDTH               (18),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk_in_clk),                     //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (33),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (45),
		.PKT_BYTE_CNT_H            (41),
		.PKT_BYTE_CNT_L            (39),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (44),
		.PKT_BURSTWRAP_L           (42),
		.PKT_TRANS_COMPRESSED_READ (34),
		.PKT_TRANS_WRITE           (36),
		.PKT_TRANS_READ            (37),
		.ST_DATA_W                 (57),
		.ST_CHANNEL_W              (18),
		.OUT_BYTE_CNT_H            (39),
		.OUT_BURSTWRAP_H           (44),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (clk_clk_in_clk),                      //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),         //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),          //          .data
		.sink0_channel         (width_adapter_002_src_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),         //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (54),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (18),
		.OUT_BYTE_CNT_H            (49),
		.OUT_BURSTWRAP_H           (53),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (clk_clk_in_clk),                          //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),                 //     sink0.valid
		.sink0_data            (width_adapter_src_data),                  //          .data
		.sink0_channel         (width_adapter_src_channel),               //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),         //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),           //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),                 //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (54),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (18),
		.OUT_BYTE_CNT_H            (49),
		.OUT_BURSTWRAP_H           (53),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_002 (
		.clk                   (clk_clk_in_clk),                          //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~clk_clk_in_reset_reset_n),                  // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk_in_clk),                             //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	system_0_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk_in_clk),                    //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket)    //           .endofpacket
	);

	system_0_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk_clk_in_clk),                         //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket)    //           .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk_in_clk),                        //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk_in_clk),                        //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk_in_clk),                        //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clk_clk_in_clk),                        //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	system_0_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (clk_clk_in_clk),                        //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk_in_clk),                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_005_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_005_src_channel),         //          .channel
		.sink_data          (width_adapter_005_src_data),            //          .data
		.sink_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_005_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_005 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_006 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_007 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_008 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_009 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_010 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_011 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_012 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_013 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_014 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_015 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_016 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_demux_005 rsp_xbar_demux_017 (
		.clk                (clk_clk_in_clk),                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk_in_clk),                        //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	system_0_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk_clk_in_clk),                        //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (68),
		.IN_PKT_BYTE_CNT_L             (66),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (71),
		.IN_PKT_BURSTWRAP_L            (69),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (50),
		.OUT_PKT_BYTE_CNT_L            (48),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (18),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk               (clk_clk_in_clk),                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid          (cmd_xbar_mux_001_src_valid),         //      sink.valid
		.in_channel        (cmd_xbar_mux_001_src_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_mux_001_src_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_mux_001_src_ready),         //          .ready
		.in_data           (cmd_xbar_mux_001_src_data),          //          .data
		.out_endofpacket   (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data          (width_adapter_src_data),             //          .data
		.out_channel       (width_adapter_src_channel),          //          .channel
		.out_valid         (width_adapter_src_valid),            //          .valid
		.out_ready         (width_adapter_src_ready),            //          .ready
		.out_startofpacket (width_adapter_src_startofpacket)     //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (50),
		.IN_PKT_BYTE_CNT_L             (48),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (53),
		.IN_PKT_BURSTWRAP_L            (51),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (68),
		.OUT_PKT_BYTE_CNT_L            (66),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (18),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk               (clk_clk_in_clk),                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid          (id_router_001_src_valid),             //      sink.valid
		.in_channel        (id_router_001_src_channel),           //          .channel
		.in_startofpacket  (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_001_src_ready),             //          .ready
		.in_data           (id_router_001_src_data),              //          .data
		.out_endofpacket   (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_001_src_data),          //          .data
		.out_channel       (width_adapter_001_src_channel),       //          .channel
		.out_valid         (width_adapter_001_src_valid),         //          .valid
		.out_ready         (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket (width_adapter_001_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (68),
		.IN_PKT_BYTE_CNT_L             (66),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (71),
		.IN_PKT_BURSTWRAP_L            (69),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (33),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (41),
		.OUT_PKT_BYTE_CNT_L            (39),
		.OUT_PKT_TRANS_COMPRESSED_READ (34),
		.OUT_ST_DATA_W                 (57),
		.ST_CHANNEL_W                  (18),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk               (clk_clk_in_clk),                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid          (cmd_xbar_mux_003_src_valid),          //      sink.valid
		.in_channel        (cmd_xbar_mux_003_src_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_mux_003_src_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_003_src_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_mux_003_src_ready),          //          .ready
		.in_data           (cmd_xbar_mux_003_src_data),           //          .data
		.out_endofpacket   (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_002_src_data),          //          .data
		.out_channel       (width_adapter_002_src_channel),       //          .channel
		.out_valid         (width_adapter_002_src_valid),         //          .valid
		.out_ready         (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket (width_adapter_002_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (33),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (41),
		.IN_PKT_BYTE_CNT_L             (39),
		.IN_PKT_TRANS_COMPRESSED_READ  (34),
		.IN_PKT_BURSTWRAP_H            (44),
		.IN_PKT_BURSTWRAP_L            (42),
		.IN_ST_DATA_W                  (57),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (68),
		.OUT_PKT_BYTE_CNT_L            (66),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (18),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_003 (
		.clk               (clk_clk_in_clk),                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid          (id_router_003_src_valid),             //      sink.valid
		.in_channel        (id_router_003_src_channel),           //          .channel
		.in_startofpacket  (id_router_003_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_003_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_003_src_ready),             //          .ready
		.in_data           (id_router_003_src_data),              //          .data
		.out_endofpacket   (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_003_src_data),          //          .data
		.out_channel       (width_adapter_003_src_channel),       //          .channel
		.out_valid         (width_adapter_003_src_valid),         //          .valid
		.out_ready         (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket (width_adapter_003_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (68),
		.IN_PKT_BYTE_CNT_L             (66),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (71),
		.IN_PKT_BURSTWRAP_L            (69),
		.IN_ST_DATA_W                  (84),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (50),
		.OUT_PKT_BYTE_CNT_L            (48),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (18),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_004 (
		.clk               (clk_clk_in_clk),                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid          (cmd_xbar_mux_004_src_valid),          //      sink.valid
		.in_channel        (cmd_xbar_mux_004_src_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_mux_004_src_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_004_src_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_mux_004_src_ready),          //          .ready
		.in_data           (cmd_xbar_mux_004_src_data),           //          .data
		.out_endofpacket   (width_adapter_004_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_004_src_data),          //          .data
		.out_channel       (width_adapter_004_src_channel),       //          .channel
		.out_valid         (width_adapter_004_src_valid),         //          .valid
		.out_ready         (width_adapter_004_src_ready),         //          .ready
		.out_startofpacket (width_adapter_004_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (50),
		.IN_PKT_BYTE_CNT_L             (48),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (53),
		.IN_PKT_BURSTWRAP_L            (51),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (68),
		.OUT_PKT_BYTE_CNT_L            (66),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_ST_DATA_W                 (84),
		.ST_CHANNEL_W                  (18),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_005 (
		.clk               (clk_clk_in_clk),                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid          (id_router_004_src_valid),             //      sink.valid
		.in_channel        (id_router_004_src_channel),           //          .channel
		.in_startofpacket  (id_router_004_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_004_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_004_src_ready),             //          .ready
		.in_data           (id_router_004_src_data),              //          .data
		.out_endofpacket   (width_adapter_005_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_005_src_data),          //          .data
		.out_channel       (width_adapter_005_src_channel),       //          .channel
		.out_valid         (width_adapter_005_src_valid),         //          .valid
		.out_ready         (width_adapter_005_src_ready),         //          .ready
		.out_startofpacket (width_adapter_005_src_startofpacket)  //          .startofpacket
	);

	system_0_irq_mapper irq_mapper (
		.clk           (clk_clk_in_clk),                 //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

endmodule
