//Componentes varios

//Banco de registros de dos salidas y una entrada
module regfile(input  wire        clk, 
               input  wire        we3,           //se�al de habilitaci�n de escritura
               input  wire [3:0]  ra1, ra2, wa3, //direcciones de regs leidos y reg a escribir
               input  wire [7:0]  wd3, 			 //dato a escribir
               output wire [7:0]  rd1, rd2);     //datos leidos

  reg [7:0] regb[0:15]; //memoria de 16 registros de 8 bits de ancho

  // El registro 0 siempre es cero
  // se leen dos reg combinacionalmente
  // y la escritura del tercero ocurre en flanco de subida del reloj
  always @(posedge clk)
    if (we3) regb[wa3] <= wd3;	
  
  assign rd1 = (ra1 != 0) ? regb[ra1] : 0;
  assign rd2 = (ra2 != 0) ? regb[ra2] : 0;
endmodule

//modulo sumador  
module sum(input  wire [9:0] a, b,
             output wire [9:0] y);

  assign y = a + b;
endmodule

//modulo de registro para modelar el PC, cambia en cada flanco de subida de reloj o de reset
module registro #(parameter WIDTH = 8)
              (input  wire             clk, reset,
               input  wire [WIDTH-1:0] d, 
               output reg  [WIDTH-1:0] q);

  always @(posedge clk, posedge reset)
    if (reset) q <= 0;
    else       q <= d;
endmodule

module registroCE #(parameter WIDTH = 8)
              (input  wire             clk, reset, enable,
               input  wire [WIDTH-1:0] d, 
               output reg  [WIDTH-1:0] q);

  always @(clk, reset, enable)
  begin
    if (reset) q <= 0;
    else 
    begin
       if ((clk==0)&(enable)) q <= d;
    end
  end
endmodule

module mux2 #(parameter WIDTH = 8)
             (input  wire [WIDTH-1:0] d0, d1, 
              input  wire             s, 
              output wire [WIDTH-1:0] y);

  assign y = s ? d1 : d0; 
endmodule

module mux4 #(parameter WIDTH = 8)
             (input  wire [WIDTH-1:0] d0, d1, d2, d3,
              input  wire [1:0]       s, 
              output wire [WIDTH-1:0] y);

  assign y = ((s[1]==0)&(s[0]==0))? d0 : ((s[1]==0)&(s[0]==1))? d1 : ((s[1]==1)&(s[0]==0))? d2 : d3;  
endmodule

module dec2(input wire           enable,
              input  wire [1:0]       s, 
              output wire y0, y1, y2, y3);
              
  assign y0 = ((s[1]==0)&(s[0]==0))? enable : 0;
  assign y1 = ((s[1]==0)&(s[0]==1))? enable : 0;
  assign y2 = ((s[1]==1)&(s[0]==0))? enable : 0;
  assign y3 = ((s[1]==1)&(s[0]==1))? enable : 0;
endmodule